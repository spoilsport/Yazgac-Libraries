* AD588 SPICE Macromodel
* Description: Reference
* Generic Desc: �5/�10Vout, 36Vin,  Zener REF, pin prog.
* Developed by: AAG / ADSC
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (04/1994)
* Copyright 1994, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include:
*
* END Notes
*
*  NODE NUMBERS
*
*       A3 OUT FORCE    =       Node 1
*       V+              =       Node 2
*       A3 OUT SENSE    =       Node 3
*       A3 +IN          =       Node 4
*       GAIN ADJ        =       Node 5
*       VHIGH           =       Node 6
*       NOISE           =       Node 7
*       VLOW            =       Node 8
*       GND SENSE +IN   =       Node 9
*       GND SENSE -IN   =       Node 10
*       VCT             =       Node 11
*       BAL ADJ         =       Node 12
*       A4 +IN          =       Node 13
*       A4 OUT SENSE    =       Node 14
*       A4 OUT FORCE    =       Node 15
*       V-              =       Node 16
*
.SUBCKT AD588 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
*
* BURIED ZENER REFERENCE CORE
*
IZ1 8 20 DC 6.848095E-3
RZ1 20 8 1E3 TC1=3E-6
ENZ 21 20 23 0 1
GZ1 8 21 2 0 1.37E-7
FZ1 8 21 POLY(4) VS1A3 VS2A3 VS1A4 VS2A4
+ (0,3.425E-5,-3.425E-5,-3.425E-5,3.425E-5)
RNR 21 7 4.2E3
*
* REFERENCE CORE VOLTAGE NOISE GENERATOR
*
VN1 22 0 DC 2
DN1 22 23 DEN1
DN2 23 24 DEN1
VN2 0 24 DC 2
*
* REFERENCE CORE AMPLIFIER A1
*
R1A1 2 30 2.122065E4
R2A1 2 31 2.122065E4
Q1A1 30 25 32 QNA1
Q2A1 31 7 33 QNA1
R3A1 32 34 2.070346E4
R4A1 33 34 2.070346E4
I1A1 34 16 DC 100E-6
*
* GAIN STAGE AND DOMINANT POLE AT 5 Hz
*
ERA1 35 0 POLY(2) 2 0 16 0 (0,0.5,0.5)
G1A1 35 36 30 31 4.712389E-5
R5A1 36 35 2.122065E9
C1A1 36 35 1.5E-11
V1A1 2 37 DC 2.5
D1A1 36 37 DX
V2A1 38 16 DC 4 
D2A1 38 36 DX
*
* OUTPUT STAGE A1
*
G2A1 35 39 36 35 1E-4
R6A1 39 35 1E4
Q3A1 2 39 40 QNA1
Q4A1 39 40 6 QNA1
R7A1 40 6 40
*
* INTERNAL RESISTOR NETWORK, GAIN AND BALANCE TRIMS
*
R1 6 25 6.3E3
R2 25 8 13.7E3
R3 5 25 150E3
IGA 5 0 DC 0
R4 6 26 10E3
R5 26 8 10E3
R6 26 12 150E3
R7 6 11 10E3
R8 11 26 150E3
R9 11 8 10E3
IBA 12 0 DC 0
ISY 2 16 DC 4.206E-3
*
* GND SENSE AMPLIFIER A2
* INPUT STAGE WITH POLE AT 3 MHz
*
EPOS 110 0 2 0 1
ENEG 120 0 16 0 1
Q1A2 41 10 43 QNA2
Q2A2 42 9 44 QNA2
R1A2 110 41 5.305096
R2A2 110 42 5.305096
C1A2 41 42 2E-8
R3A2 43 45 0.133096
R4A2 44 45 0.133096
I1A2 45 120 DC 1E-2
*
* GAIN STAGE AND DOMINANT POLE AT 3.1623 Hz
*
ERA2 46 0 POLY(2) 2 0 16 0 (0,0.5,0.5)
G1A2 46 47 41 42 1.88498E-1
R5A2 47 46 1.67763E6
C2A2 47 46 3E-8
V1A2 110 48 DC 2.2
D1A2 47 48 DX
V2A2 49 120 DC 2.2
D2A2 49 47 DX
*
* OUTPUT STAGE A2
*
E1A2 50 46 47 46 1
Q3A2 16 50 8 QPA2
*
* OUTPUT AMPLIFIER A3
*
R1A3 3 51 1E6
R2A3 51 4 1E6
R3A3 2 52 530.5096
R4A3 2 53 530.5096
Q1A3 52 3 54 QNA3
Q2A3 53 58 55 QNA3
R5A3 54 56 13.3096
R6A3 55 56 13.3096
EOSA3 57 4 POLY(1) 67 62 (100E-6,1)
ENA3 58 57 60 0 1
I1A3 56 16 DC 100E-6
*
* A3 INPUT VOLTAGE NOISE GENERATOR
*
VN1A3 59 0 DC 2
DN1A3 59 60 DEN2
DN2A3 60 61 DEN2
VN2A3 0 61 DC 2
*
* GAIN STAGE AND DOMINANT POLE AT 3.1623 Hz
*
ERA3 62 0 POLY(2) 2 0 16 0 (0,0.5,0.5)
G1A3 62 63 52 53 1.88498E-3
R7A3 63 62 1.67763E8
C1A3 63 62 3E-10
V1A3 2 64 DC 3.5
D1A3 63 64 DX
V2A3 65 16 DC 3.5
D2A3 65 63 DX
*
* COMMON-MODE REJECTION STAGE AND ZERO AT 2 kHz
*
ECMA3 66 62 51 62 10
RCM1A3 66 67 1E6
CCMA3 66 67 7.9577E-11
RCM2A3 67 62 1
*
* POLE AT 2.5 MHz
*
G2A3 62 68 63 62 1E-6
R8A3 68 62 1E6
C2A3 68 62 6.3662E-14
*
* A3 OUTPUT STAGE
*
DSC1A3 68 69 DX
VSC1A3 69 71 DC 4.4
DSC2A3 70 68 DX
VSC2A3 71 70 DC 4.4
FSYA3 2 16 POLY(2) VSY1A3 VSY2A3 (0,1,1)
GSYA3 62 74 71 68 5E-3
DSY1A3 74 75 DX
VSY1A3 75 62 DC 0
DSY2A3 76 74 DX
VSY2A3 62 76 DC 0
GO1A3 71 2 2 68 5E-3
RO1A3 2 71 200
GO2A3 16 71 68 16 5E-3
RO2A3 16 71 200
VOA3 72 71 DC 0
FA3 62 73 VOA3 1
DS1A3 73 103 DX
VS1A3 103 62 DC 0
DS2A3 104 73 DX
VS2A3 62 104 DC 0
L1A3 72 1 1E-7
*
* OUTPUT AMPLIFIER A4
*
R1A4 14 77 1E6
R2A4 77 13 1E6
R3A4 2 78 530.5096
R4A4 2 79 530.5096
Q1A4 78 14 80 QNA3
Q2A4 79 84 81 QNA3
R5A4 80 82 13.3096
R6A4 81 82 13.3096
EOSA4 83 13 POLY(1) 93 88 (100E-6,1)
ENA4 84 83 86 0 1
I1A4 82 16 DC 100E-6
*
* A4 INPUT VOLTAGE NOISE GENERATOR
*
VN1A4 85 0 DC 2
DN1A4 85 86 DEN2
DN2A4 86 87 DEN2
VN2A4 0 87 DC 2
*
* GAIN STAGE AND DOMINANT POLE AT 3.1623 Hz
*
ERA4 88 0 POLY(2) 2 0 16 0 (0,0.5,0.5)
G1A4 88 89 78 79 1.88498E-3
R7A4 89 88 1.67763E8
C1A4 89 88 3E-10
V1A4 2 90 DC 3.5
D1A4 89 90 DX
V2A4 91 16 DC 3.5
D2A4 91 89 DX
*
* COMMON-MODE REJECTION STAGE AND ZERO AT 2 kHz
*
ECMA4 92 88 77 88 10
RCM1A4 92 93 1E6
CCMA4 92 93 7.9577E-11
RCM2A4 93 88 1
*
* POLE AT 2.5 MHz
*
G2A4 88 94 89 88 1E-6
R8A4 94 88 1E6
C2A4 94 88 6.3662E-14
*
* A4 OUTPUT STAGE
*
DSC1A4 94 95 DX
VSC1A4 95 97 DC 4.4
DSC2A4 96 94 DX
VSC2A4 97 96 DC 4.4
FSYA4 2 16 POLY(2) VSY1A4 VSY2A4 (0,1,1)
GSYA4 88 100 97 94 5E-3
DSY1A4 100 101 DX
VSY1A4 101 88 DC 0
DSY2A4 102 100 DX
VSY2A4 88 102 DC 0
GO1A4 97 2 2 94 5E-3
RO1A4 2 97 200
GO2A4 16 97 94 16 5E-3
RO2A4 16 97 200
VOA4 98 97 DC 0
FA4 88 99 VOA4 1
DS1A4 99 105 DX
VS1A4 105 88 DC 0
DS2A4 106 99 DX
VS2A4 88 106 DC 0
L1A4 98 15 1E-7
*
.MODEL QNA1 NPN(IS=1E-15 BF=1E3)
.MODEL QNA2 NPN(IS=1E-15 BF=2.5E5)
.MODEL QNA3 NPN(IS=1E-15 BF=2.5E3)
.MODEL QPA2 PNP(IS=1E-15 BF=1E3)
.MODEL DX D(IS=1E-15)
.MODEL DEN1 D(IS=1E-12 RS=2.87035E+05 AF=1 KF=1.15709E-15)
.MODEL DEN2 D(IS=1E-12 RS=1.903E+05 AF=1 KF=2.200E-16)
*
.ENDS AD588






